module memory #(parameter C=256, W=32) (input [W-1:0] data,input [7:0] ad,input WE,clk, output reg [W-1:0] RD);

reg [W-1:0] mem [C-1:0];

initial begin
//mem[8'h00]=17'b01100000100000001;
//mem[8'h01]=17'b00000101100101000;

mem[8'h00]=17'b00010101000000000;
mem[8'h01]=17'b01110000100001100;
mem[8'h02]=17'b01110000100001100;
mem[8'h03]=17'b01110000100001110;
mem[8'h04]=17'b00000001000101000;
mem[8'h05]=17'b01110000100001110;
mem[8'h06]=17'b00000001000101000;
mem[8'h07]=17'b01110000100001111;
mem[8'h08]=17'b00000001000101000;
mem[8'h09]=17'b01110000100010000;
mem[8'h0A]=17'b00000001000101000;
mem[8'h0B]=17'b01000001000010001;

mem[8'h0C]=17'b00000000000000011;
mem[8'h0D]=17'b00000000000000111;
mem[8'h0E]=17'b00000000000001001;
mem[8'h0F]=17'b00000000000000001;
mem[8'h10]=17'b00000000000001110;



end

always @(posedge clk)
	if(WE)
		mem[ad]<=data;
		

always @(*)
	RD=mem[ad];
	
endmodule